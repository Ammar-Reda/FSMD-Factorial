library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;

entity mux_2_1_13bit is
    port (s: in std_logic;
            a, b: in std_logic_vector(12 downto 0);
            y: out std_logic_vector(12 downto 0));
end entity mux_2_1_13bit;

architecture rtl of mux_2_1_13bit is
begin

y <= a when s = '0' else b;

end architecture rtl;
